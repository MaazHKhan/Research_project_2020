when s0 => -- intialisation state
	x <= -524288;
	state <= s1;
	report "In state 0";